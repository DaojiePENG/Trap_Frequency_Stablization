`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: SUSTech
// Engineer: Daojie.PENG@outlook.com
// 
// Create Date: 2023年3月20日04:14:22
// Design Name: 
// Module Name: Full_Ahead_2Adder
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: carray ahead adder 
//            it has 0 pipeline stage
// Dependencies: full_ahead_adder
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// Reference： https://blog.csdn.net/qq_26707507/article/details/106146619
//////////////////////////////////////////////////////////////////////////////////

module Full_Ahead_2Adder #(
    parameter Width = 64,// width of the ahead adder, it can be 2, 4, 8, 16, 32, 64.
    parameter Stage = 0)(
    input  wire             i_clkp  ,
    input  wire             i_rstn  ,
    input  wire             i_c     , // 前一级进位
    input  wire [Width-1:0] i_a     , // 被加数
    input  wire [Width-1:0] i_b     , // 加数

    output wire [Width-1:0] o_d     , // 和
    output wire             o_c     , // 进位
    output wire             o_gm    , // generater of MSB
    output wire             o_pm      // propagater of MSB
    );
/*
carray look ahead adder
*/
wire [Width-1:0] g_wire, p_wire, d_wire;
wire [Width:0] c_wire;
assign c_wire[0]=i_c;

generate
    genvar i;
    for (i = 0; i < Width; i = i + 1)
        begin: ahead_adder4_gene
            full_adder1 adder(
                .i_c    (c_wire [i] ),
                .i_a    (i_a    [i] ),
                .i_b    (i_b    [i] ),

                .o_d    (d_wire [i] ),
                .o_g    (g_wire [i] ),
                .o_p    (p_wire [i] ) 
                );
        end
endgenerate
wire gm_wire, pm_wire;
generate// generate different encoders based on Width
    if (Width==2)
        begin
            carray_ahead_encoder2 encoder2(// encoder for carray ahead adder.
                .i_c    (i_c            ),
                .i_g    (g_wire         ),
                .i_p    (p_wire         ),

                .o_c    (c_wire[Width:1]),
                .o_gm   (gm_wire        ),
                .o_pm   (pm_wire        )         
                );
        end
    else if (Width==4)
        begin
            carray_ahead_encoder4 encoder4(// encoder for carray ahead adder.
                .i_c    (i_c            ),
                .i_g    (g_wire         ),
                .i_p    (p_wire         ),

                .o_c    (c_wire[Width:1]),
                .o_gm   (gm_wire        ),
                .o_pm   (pm_wire        )         
                );
        end
    else if (Width==8)
        begin
            carray_ahead_encoder8 encoder8(// encoder for carray ahead adder.
                .i_c    (i_c            ),
                .i_g    (g_wire         ),
                .i_p    (p_wire         ),

                .o_c    (c_wire[Width:1]),
                .o_gm   (gm_wire        ),
                .o_pm   (pm_wire        )         
                );
        end
    else if (Width==16)
        begin
            carray_ahead_encoder16 encoder16(// encoder for carray ahead adder.
                .i_c    (i_c            ),
                .i_g    (g_wire         ),
                .i_p    (p_wire         ),

                .o_c    (c_wire[Width:1]),
                .o_gm   (gm_wire        ),
                .o_pm   (pm_wire        )         
                );
        end
    else if (Width==32)
        begin
            carray_ahead_encoder32 encoder32(// encoder for carray ahead adder.
                .i_c    (i_c            ),
                .i_g    (g_wire         ),
                .i_p    (p_wire         ),

                .o_c    (c_wire[Width:1]),
                .o_gm   (gm_wire        ),
                .o_pm   (pm_wire        )         
                );
        end
    else if (Width==64)
        begin
            carray_ahead_encoder64 encoder64(// encoder for carray ahead adder.
                .i_c    (i_c            ),
                .i_g    (g_wire         ),
                .i_p    (p_wire         ),

                .o_c    (c_wire[Width:1]),
                .o_gm   (gm_wire        ),
                .o_pm   (pm_wire        )         
                );
        end
endgenerate

pipelineto  #(.Width(Width+3),.Stage(Stage)) lineto_output(// choose output pipeline
  .i_clkp(i_clkp), .i_rstn(i_rstn),
  .i_a({d_wire, c_wire[Width],  gm_wire,    pm_wire }),
  .o_a({o_d,    o_c,            o_gm,       o_pm    })
  );
/*
assign o_d=d_wire;
assign o_c=c_wire[Width];
assign o_gm=gm_wire;
assign o_pm=pm_wire;
*/
endmodule


/**/

//////////////////////////////////////////////////////////////////////////////////
// Company: SUSTech
// Engineer: Daojie.PENG@qq.com
// 
// Create Date: 2022/09/15 20:46:40
// Design Name: full adder1 
// Module Name: full_adder1 
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: full adder for carray lookahead adder encoding 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module full_adder1(// adder for carray ahead adder
    input  wire i_c     , // carry in
    input  wire i_a     , // augend
    input  wire i_b     , // addend

    output wire o_d     , // sum out
    output wire o_g     , // generater
    output wire o_p       // propagter
    );
    assign o_d = i_a ^ i_b ^ i_c;
    assign o_g = i_a & i_b; // 
    assign o_p = i_a ^ i_b; // work with carray in
endmodule


//////////////////////////////////////////////////////////////////////////////////
// Company: SUSTech
// Engineer: Daojie.PENG@qq.com
// 
// Create Date: 2022/09/15 20:46:40
// Design Name: carray_ahead_encoder
// Module Name: carray_ahead_encoder 
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: encoder for carray lookahead adder encoding 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

//2位CLA部件
module carray_ahead_encoder2(// use genearter and propagater to get the look-ahead carray of each bit
    input           i_c     ,
    input [1:0]     i_g     ,
    input [1:0]     i_p     ,

    output [2:1]    o_c     ,
    output          o_gm    ,
    output          o_pm     
    );
assign o_c[1]=i_g[0] | i_p[0]&i_c;
assign o_c[2]=i_g[1] | i_p[1]&i_g[0] | i_p[1]&i_p[0]&i_c;

assign o_gm=i_g[1] | i_p[1]&i_g[0] ;// generater of MSB
assign o_pm=i_p[1]&i_p[0];// propagater of MSB
endmodule


//4位CLA部件
module carray_ahead_encoder4(// use genearter and propagater to get the look-ahead carray of each bit
    input           i_c     ,
    input [3:0]     i_g     ,
    input [3:0]     i_p     ,

    output [4:1]    o_c     ,
    output          o_gm    ,
    output          o_pm    
    );
assign o_c[1]=i_g[0] | i_p[0]&i_c;
assign o_c[2]=i_g[1] | i_p[1]&i_g[0] | i_p[1]&i_p[0]&i_c;
assign o_c[3]=i_g[2] | i_p[2]&i_g[1] | i_p[2]&i_p[1]&i_g[0] | i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[4]=i_g[3] | i_p[3]&i_g[2] | i_p[3]&i_p[2]&i_g[1] | i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;

assign o_gm=i_g[3] | i_p[3]&i_g[2] | i_p[3]&i_p[2]&i_g[1] | i_p[3]&i_p[2]&i_p[1]&i_g[0];// generater of MSB
assign o_pm=i_p[3]&i_p[2]&i_p[1]&i_p[0];// propagater of MSB
endmodule

/*
module carray_ahead_encoder4_1(// use genearter and propagater to get the look-ahead carray of each bit
    input           i_c     ,
    input [3:0]     i_g     ,
    input [3:0]     i_p     ,

    output [4:1]    o_c     ,
    output          o_gm    ,
    output          o_pm    
    );
assign o_c[1]=i_g[0] | i_p[0]&i_c;
assign o_c[2]=i_g[1] | i_p[1]&o_c[1];
assign o_c[3]=i_g[2] | i_p[2]&o_c[2];
assign o_c[4]=i_g[3] | i_p[3]&o_c[3];

assign o_gm=i_g[3] | i_p[3]&i_g[2] | i_p[3]&i_p[2]&i_g[1] | i_p[3]&i_p[2]&i_p[1]&i_g[0];// generater of MSB
assign o_pm=i_p[3]&i_p[2]&i_p[1]&i_p[0];// propagater of MSB
endmodule
*/

//8位CLA部件
module carray_ahead_encoder8(// use genearter and propagater to get the look-ahead carray of each bit
    input           i_c     ,
    input [7:0]     i_g     ,
    input [7:0]     i_p     ,

    output [8:1]    o_c     ,
    output          o_gm    ,
    output          o_pm    
    );
assign o_c[1]=i_g[0] | i_p[0]&i_c;
assign o_c[2]=i_g[1] | i_p[1]&i_g[0] | i_p[1]&i_p[0]&i_c;
assign o_c[3]=i_g[2] | i_p[2]&i_g[1] | i_p[2]&i_p[1]&i_g[0] | i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[4]=i_g[3] | i_p[3]&i_g[2] | i_p[3]&i_p[2]&i_g[1] | i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;

// 要继续拓展的规律为每次前面 | 上生成子i_g，然后上一级的所有 & 上传输子i_p; 各级以此类推
assign o_c[5]=i_g[4] | i_p[4]&i_g[3] | i_p[4]&i_p[3]&i_g[2] | i_p[4]&i_p[3]&i_p[2]&i_g[1] | i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[6]=i_g[5] | i_p[5]&i_g[4] | i_p[5]&i_p[4]&i_g[3] | i_p[5]&i_p[4]&i_p[3]&i_g[2] | i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_g[1] | i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[7]=i_g[6] | i_p[6]&i_g[5] | i_p[6]&i_p[5]&i_g[4] | i_p[6]&i_p[5]&i_p[4]&i_g[3] | i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_g[2] | i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_g[1] | i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[8]=i_g[7] | i_p[7]&i_g[6] | i_p[7]&i_p[6]&i_g[5] | i_p[7]&i_p[6]&i_p[5]&i_g[4] | i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_g[3] | i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_g[2] | i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_g[1] | i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;

assign o_gm=i_g[7] | i_p[7]&i_g[6] | i_p[7]&i_p[6]&i_g[5] | i_p[7]&i_p[6]&i_p[5]&i_g[4] | i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_g[3] | i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_g[2] | i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_g[1] | i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_g[0];// generater of MSB
assign o_pm=i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0];// propagater of MSB
endmodule

//16位CLA部件
module carray_ahead_encoder16(// use genearter and propagater to get the look-ahead carray of each bit
    input           i_c     ,
    input  [15:0]   i_g     ,
    input  [15:0]   i_p     ,

    output [16:1]   o_c     ,
    output          o_gm    ,
    output          o_pm    
    );
assign o_c[1]=i_g[0] | i_p[0]&i_c;
assign o_c[2]=i_g[1] | i_p[1]&i_g[0] | i_p[1]&i_p[0]&i_c;
assign o_c[3]=i_g[2] | i_p[2]&i_g[1] | i_p[2]&i_p[1]&i_g[0] | i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[4]=i_g[3] | i_p[3]&i_g[2] | i_p[3]&i_p[2]&i_g[1] | i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;

// 要继续拓展的规律为每次前面 | 上生成子i_g，然后上一级的所有 & 上传输子i_p; 各级以此类推
assign o_c[ 5]=i_g[4] | i_p[4]&i_g[3] | i_p[4]&i_p[3]&i_g[2] | i_p[4]&i_p[3]&i_p[2]&i_g[1] | i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[ 6]=i_g[5] | i_p[5]&i_g[4] | i_p[5]&i_p[4]&i_g[3] | i_p[5]&i_p[4]&i_p[3]&i_g[2] | i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_g[1] | i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[ 7]=i_g[6] | i_p[6]&i_g[5] | i_p[6]&i_p[5]&i_g[4] | i_p[6]&i_p[5]&i_p[4]&i_g[3] | i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_g[2] | i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_g[1] | i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[ 8]=i_g[7] | i_p[7]&i_g[6] | i_p[7]&i_p[6]&i_g[5] | i_p[7]&i_p[6]&i_p[5]&i_g[4] | i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_g[3] | i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_g[2] | i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_g[1] | i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[ 9]=i_g[8] | i_p[8]&i_g[7] | i_p[8]&i_p[7]&i_g[6] | i_p[8]&i_p[7]&i_p[6]&i_g[5] | i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_g[4] | i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_g[3] | i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_g[2] | i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_g[1] | i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[10]=i_g[9] | i_p[9]&i_g[8] | i_p[9]&i_p[8]&i_g[7] | i_p[9]&i_p[8]&i_p[7]&i_g[6] | i_p[9]&i_p[8]&i_p[7]&i_p[6]&i_g[5] | i_p[9]&i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_g[4] | i_p[9]&i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_g[3] | i_p[9]&i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_g[2] | i_p[9]&i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_g[1] | i_p[9]&i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[9]&i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[11]=i_g[10] | i_p[10]&i_g[ 9] | i_p[10]&i_p[ 9]&i_g[ 8] | i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[12]=i_g[11] | i_p[11]&i_g[10] | i_p[11]&i_p[10]&i_g[ 9] | i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[13]=i_g[12] | i_p[12]&i_g[11] | i_p[12]&i_p[11]&i_g[10] | i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[14]=i_g[13] | i_p[13]&i_g[12] | i_p[13]&i_p[12]&i_g[11] | i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[15]=i_g[14] | i_p[14]&i_g[13] | i_p[14]&i_p[13]&i_g[12] | i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[16]=i_g[15] | i_p[15]&i_g[14] | i_p[15]&i_p[14]&i_g[13] | i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;


assign o_gm=i_g[15] | i_p[15]&i_g[14] | i_p[15]&i_p[14]&i_g[13] | i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0];// generater of MSB
assign o_pm=i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[9]&i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0];// propagater of MSB
endmodule

//32位CLA部件
module carray_ahead_encoder32(// use genearter and propagater to get the look-ahead carray of each bit
    input           i_c     ,
    input  [31:0]   i_g     ,
    input  [31:0]   i_p     ,

    output [32:1]   o_c     ,
    output          o_gm    ,
    output          o_pm    
    );
assign o_c[1]=i_g[0] | i_p[0]&i_c;
assign o_c[2]=i_g[1] | i_p[1]&i_g[0] | i_p[1]&i_p[0]&i_c;
assign o_c[3]=i_g[2] | i_p[2]&i_g[1] | i_p[2]&i_p[1]&i_g[0] | i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[4]=i_g[3] | i_p[3]&i_g[2] | i_p[3]&i_p[2]&i_g[1] | i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;

// 要继续拓展的规律为每次前面 | 上生成子i_g，然后上一级的所有 & 上传输子i_p; 各级以此类推
assign o_c[ 5]=i_g[4] | i_p[4]&i_g[3] | i_p[4]&i_p[3]&i_g[2] | i_p[4]&i_p[3]&i_p[2]&i_g[1] | i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[ 6]=i_g[5] | i_p[5]&i_g[4] | i_p[5]&i_p[4]&i_g[3] | i_p[5]&i_p[4]&i_p[3]&i_g[2] | i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_g[1] | i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[ 7]=i_g[6] | i_p[6]&i_g[5] | i_p[6]&i_p[5]&i_g[4] | i_p[6]&i_p[5]&i_p[4]&i_g[3] | i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_g[2] | i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_g[1] | i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[ 8]=i_g[7] | i_p[7]&i_g[6] | i_p[7]&i_p[6]&i_g[5] | i_p[7]&i_p[6]&i_p[5]&i_g[4] | i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_g[3] | i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_g[2] | i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_g[1] | i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[ 9]=i_g[8] | i_p[8]&i_g[7] | i_p[8]&i_p[7]&i_g[6] | i_p[8]&i_p[7]&i_p[6]&i_g[5] | i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_g[4] | i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_g[3] | i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_g[2] | i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_g[1] | i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[10]=i_g[9] | i_p[9]&i_g[8] | i_p[9]&i_p[8]&i_g[7] | i_p[9]&i_p[8]&i_p[7]&i_g[6] | i_p[9]&i_p[8]&i_p[7]&i_p[6]&i_g[5] | i_p[9]&i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_g[4] | i_p[9]&i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_g[3] | i_p[9]&i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_g[2] | i_p[9]&i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_g[1] | i_p[9]&i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[9]&i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[11]=i_g[10] | i_p[10]&i_g[ 9] | i_p[10]&i_p[ 9]&i_g[ 8] | i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[12]=i_g[11] | i_p[11]&i_g[10] | i_p[11]&i_p[10]&i_g[ 9] | i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[13]=i_g[12] | i_p[12]&i_g[11] | i_p[12]&i_p[11]&i_g[10] | i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[14]=i_g[13] | i_p[13]&i_g[12] | i_p[13]&i_p[12]&i_g[11] | i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[15]=i_g[14] | i_p[14]&i_g[13] | i_p[14]&i_p[13]&i_g[12] | i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[16]=i_g[15] | i_p[15]&i_g[14] | i_p[15]&i_p[14]&i_g[13] | i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;

assign o_c[17]=i_g[16] | i_p[16]&i_g[15] | i_p[16]&i_p[15]&i_g[14] | i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[18]=i_g[17] | i_p[17]&i_g[16] | i_p[17]&i_p[16]&i_g[15] | i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[19]=i_g[18] | i_p[18]&i_g[17] | i_p[18]&i_p[17]&i_g[16] | i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[20]=i_g[19] | i_p[19]&i_g[18] | i_p[19]&i_p[18]&i_g[17] | i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[21]=i_g[20] | i_p[20]&i_g[19] | i_p[20]&i_p[19]&i_g[18] | i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[22]=i_g[21] | i_p[21]&i_g[20] | i_p[21]&i_p[20]&i_g[19] | i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[23]=i_g[22] | i_p[22]&i_g[21] | i_p[22]&i_p[21]&i_g[20] | i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[24]=i_g[23] | i_p[23]&i_g[22] | i_p[23]&i_p[22]&i_g[21] | i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[25]=i_g[24] | i_p[24]&i_g[23] | i_p[24]&i_p[23]&i_g[22] | i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[26]=i_g[25] | i_p[25]&i_g[24] | i_p[25]&i_p[24]&i_g[23] | i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[27]=i_g[26] | i_p[26]&i_g[25] | i_p[26]&i_p[25]&i_g[24] | i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[28]=i_g[27] | i_p[27]&i_g[26] | i_p[27]&i_p[26]&i_g[25] | i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[29]=i_g[28] | i_p[28]&i_g[27] | i_p[28]&i_p[27]&i_g[26] | i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[30]=i_g[29] | i_p[29]&i_g[28] | i_p[29]&i_p[28]&i_g[27] | i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[31]=i_g[30] | i_p[30]&i_g[29] | i_p[30]&i_p[29]&i_g[28] | i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[32]=i_g[31] | i_p[31]&i_g[30] | i_p[31]&i_p[30]&i_g[29] | i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;


assign o_gm=i_g[31] | i_p[31]&i_g[30] | i_p[31]&i_p[30]&i_g[29] | i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0];
assign o_pm=i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[9]&i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0];// propagater of MSB
endmodule

//64位CLA部件
module carray_ahead_encoder64(// use genearter and propagater to get the look-ahead carray of each bit
    input           i_c     ,
    input  [63:0]   i_g     ,
    input  [63:0]   i_p     ,

    output [64:1]   o_c     ,
    output          o_gm    ,
    output          o_pm    
    );
assign o_c[1]=i_g[0] | i_p[0]&i_c;
assign o_c[2]=i_g[1] | i_p[1]&i_g[0] | i_p[1]&i_p[0]&i_c;
assign o_c[3]=i_g[2] | i_p[2]&i_g[1] | i_p[2]&i_p[1]&i_g[0] | i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[4]=i_g[3] | i_p[3]&i_g[2] | i_p[3]&i_p[2]&i_g[1] | i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;

// 要继续拓展的规律为每次前面 | 上生成子i_g，然后上一级的所有 & 上传输子i_p; 各级以此类推
assign o_c[ 5]=i_g[4] | i_p[4]&i_g[3] | i_p[4]&i_p[3]&i_g[2] | i_p[4]&i_p[3]&i_p[2]&i_g[1] | i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[ 6]=i_g[5] | i_p[5]&i_g[4] | i_p[5]&i_p[4]&i_g[3] | i_p[5]&i_p[4]&i_p[3]&i_g[2] | i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_g[1] | i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[ 7]=i_g[6] | i_p[6]&i_g[5] | i_p[6]&i_p[5]&i_g[4] | i_p[6]&i_p[5]&i_p[4]&i_g[3] | i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_g[2] | i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_g[1] | i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[ 8]=i_g[7] | i_p[7]&i_g[6] | i_p[7]&i_p[6]&i_g[5] | i_p[7]&i_p[6]&i_p[5]&i_g[4] | i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_g[3] | i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_g[2] | i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_g[1] | i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[ 9]=i_g[8] | i_p[8]&i_g[7] | i_p[8]&i_p[7]&i_g[6] | i_p[8]&i_p[7]&i_p[6]&i_g[5] | i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_g[4] | i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_g[3] | i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_g[2] | i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_g[1] | i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[10]=i_g[9] | i_p[9]&i_g[8] | i_p[9]&i_p[8]&i_g[7] | i_p[9]&i_p[8]&i_p[7]&i_g[6] | i_p[9]&i_p[8]&i_p[7]&i_p[6]&i_g[5] | i_p[9]&i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_g[4] | i_p[9]&i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_g[3] | i_p[9]&i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_g[2] | i_p[9]&i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_g[1] | i_p[9]&i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_g[0] | i_p[9]&i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0]&i_c;
assign o_c[11]=i_g[10] | i_p[10]&i_g[ 9] | i_p[10]&i_p[ 9]&i_g[ 8] | i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[12]=i_g[11] | i_p[11]&i_g[10] | i_p[11]&i_p[10]&i_g[ 9] | i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[13]=i_g[12] | i_p[12]&i_g[11] | i_p[12]&i_p[11]&i_g[10] | i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[14]=i_g[13] | i_p[13]&i_g[12] | i_p[13]&i_p[12]&i_g[11] | i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[15]=i_g[14] | i_p[14]&i_g[13] | i_p[14]&i_p[13]&i_g[12] | i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[16]=i_g[15] | i_p[15]&i_g[14] | i_p[15]&i_p[14]&i_g[13] | i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;

assign o_c[17]=i_g[16] | i_p[16]&i_g[15] | i_p[16]&i_p[15]&i_g[14] | i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[18]=i_g[17] | i_p[17]&i_g[16] | i_p[17]&i_p[16]&i_g[15] | i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[19]=i_g[18] | i_p[18]&i_g[17] | i_p[18]&i_p[17]&i_g[16] | i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[20]=i_g[19] | i_p[19]&i_g[18] | i_p[19]&i_p[18]&i_g[17] | i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[21]=i_g[20] | i_p[20]&i_g[19] | i_p[20]&i_p[19]&i_g[18] | i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[22]=i_g[21] | i_p[21]&i_g[20] | i_p[21]&i_p[20]&i_g[19] | i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[23]=i_g[22] | i_p[22]&i_g[21] | i_p[22]&i_p[21]&i_g[20] | i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[24]=i_g[23] | i_p[23]&i_g[22] | i_p[23]&i_p[22]&i_g[21] | i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[25]=i_g[24] | i_p[24]&i_g[23] | i_p[24]&i_p[23]&i_g[22] | i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[26]=i_g[25] | i_p[25]&i_g[24] | i_p[25]&i_p[24]&i_g[23] | i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[27]=i_g[26] | i_p[26]&i_g[25] | i_p[26]&i_p[25]&i_g[24] | i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[28]=i_g[27] | i_p[27]&i_g[26] | i_p[27]&i_p[26]&i_g[25] | i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[29]=i_g[28] | i_p[28]&i_g[27] | i_p[28]&i_p[27]&i_g[26] | i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[30]=i_g[29] | i_p[29]&i_g[28] | i_p[29]&i_p[28]&i_g[27] | i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[31]=i_g[30] | i_p[30]&i_g[29] | i_p[30]&i_p[29]&i_g[28] | i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[32]=i_g[31] | i_p[31]&i_g[30] | i_p[31]&i_p[30]&i_g[29] | i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;


assign o_c[33]=i_g[32] | i_p[32]&i_g[31] | i_p[32]&i_p[31]&i_g[30] | i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[34]=i_g[33] | i_p[33]&i_g[32] | i_p[33]&i_p[32]&i_g[31] | i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[35]=i_g[34] | i_p[34]&i_g[33] | i_p[34]&i_p[33]&i_g[32] | i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[36]=i_g[35] | i_p[35]&i_g[34] | i_p[35]&i_p[34]&i_g[33] | i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[37]=i_g[36] | i_p[36]&i_g[35] | i_p[36]&i_p[35]&i_g[34] | i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[38]=i_g[37] | i_p[37]&i_g[36] | i_p[37]&i_p[36]&i_g[35] | i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[39]=i_g[38] | i_p[38]&i_g[37] | i_p[38]&i_p[37]&i_g[36] | i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[40]=i_g[39] | i_p[39]&i_g[38] | i_p[39]&i_p[38]&i_g[37] | i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;

assign o_c[41]=i_g[40] | i_p[40]&i_g[39] | i_p[40]&i_p[39]&i_g[38] | i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[42]=i_g[41] | i_p[41]&i_g[40] | i_p[41]&i_p[40]&i_g[39] | i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[43]=i_g[42] | i_p[42]&i_g[41] | i_p[42]&i_p[41]&i_g[40] | i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[44]=i_g[43] | i_p[43]&i_g[42] | i_p[43]&i_p[42]&i_g[41] | i_p[43]&i_p[42]&i_p[41]&i_g[40] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[45]=i_g[44] | i_p[44]&i_g[43] | i_p[44]&i_p[43]&i_g[42] | i_p[44]&i_p[43]&i_p[42]&i_g[41] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_g[40] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[46]=i_g[45] | i_p[45]&i_g[44] | i_p[45]&i_p[44]&i_g[43] | i_p[45]&i_p[44]&i_p[43]&i_g[42] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_g[41] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_g[40] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[47]=i_g[46] | i_p[46]&i_g[45] | i_p[46]&i_p[45]&i_g[44] | i_p[46]&i_p[45]&i_p[44]&i_g[43] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_g[42] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_g[41] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_g[40] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[48]=i_g[47] | i_p[47]&i_g[46] | i_p[47]&i_p[46]&i_g[45] | i_p[47]&i_p[46]&i_p[45]&i_g[44] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_g[43] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_g[42] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_g[41] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_g[40] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;

assign o_c[49]=i_g[48] | i_p[48]&i_g[47] | i_p[48]&i_p[47]&i_g[46] | i_p[48]&i_p[47]&i_p[46]&i_g[45] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_g[44] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_g[43] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_g[42] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_g[41] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_g[40] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[50]=i_g[49] | i_p[49]&i_g[48] | i_p[49]&i_p[48]&i_g[47] | i_p[49]&i_p[48]&i_p[47]&i_g[46] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_g[45] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_g[44] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_g[43] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_g[42] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_g[41] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_g[40] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[51]=i_g[50] | i_p[50]&i_g[49] | i_p[50]&i_p[49]&i_g[48] | i_p[50]&i_p[49]&i_p[48]&i_g[47] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_g[46] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_g[45] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_g[44] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_g[43] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_g[42] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_g[41] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_g[40] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[52]=i_g[51] | i_p[51]&i_g[50] | i_p[51]&i_p[50]&i_g[49] | i_p[51]&i_p[50]&i_p[49]&i_g[48] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_g[47] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_g[46] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_g[45] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_g[44] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_g[43] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_g[42] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_g[41] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_g[40] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[53]=i_g[52] | i_p[52]&i_g[51] | i_p[52]&i_p[51]&i_g[50] | i_p[52]&i_p[51]&i_p[50]&i_g[49] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_g[48] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_g[47] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_g[46] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_g[45] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_g[44] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_g[43] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_g[42] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_g[41] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_g[40] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[54]=i_g[53] | i_p[53]&i_g[52] | i_p[53]&i_p[52]&i_g[51] | i_p[53]&i_p[52]&i_p[51]&i_g[50] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_g[49] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_g[48] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_g[47] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_g[46] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_g[45] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_g[44] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_g[43] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_g[42] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_g[41] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_g[40] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[55]=i_g[54] | i_p[54]&i_g[53] | i_p[54]&i_p[53]&i_g[52] | i_p[54]&i_p[53]&i_p[52]&i_g[51] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_g[50] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_g[49] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_g[48] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_g[47] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_g[46] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_g[45] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_g[44] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_g[43] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_g[42] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_g[41] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_g[40] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[56]=i_g[55] | i_p[55]&i_g[54] | i_p[55]&i_p[54]&i_g[53] | i_p[55]&i_p[54]&i_p[53]&i_g[52] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_g[51] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_g[50] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_g[49] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_g[48] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_g[47] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_g[46] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_g[45] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_g[44] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_g[43] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_g[42] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_g[41] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_g[40] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;

assign o_c[57]=i_g[56] | i_p[56]&i_g[55] | i_p[56]&i_p[55]&i_g[54] | i_p[56]&i_p[55]&i_p[54]&i_g[53] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_g[52] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_g[51] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_g[50] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_g[49] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_g[48] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_g[47] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_g[46] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_g[45] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_g[44] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_g[43] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_g[42] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_g[41] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_g[40] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[58]=i_g[57] | i_p[57]&i_g[56] | i_p[57]&i_p[56]&i_g[55] | i_p[57]&i_p[56]&i_p[55]&i_g[54] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_g[53] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_g[52] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_g[51] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_g[50] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_g[49] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_g[48] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_g[47] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_g[46] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_g[45] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_g[44] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_g[43] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_g[42] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_g[41] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_g[40] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[59]=i_g[58] | i_p[58]&i_g[57] | i_p[58]&i_p[57]&i_g[56] | i_p[58]&i_p[57]&i_p[56]&i_g[55] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_g[54] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_g[53] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_g[52] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_g[51] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_g[50] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_g[49] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_g[48] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_g[47] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_g[46] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_g[45] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_g[44] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_g[43] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_g[42] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_g[41] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_g[40] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[60]=i_g[59] | i_p[59]&i_g[58] | i_p[59]&i_p[58]&i_g[57] | i_p[59]&i_p[58]&i_p[57]&i_g[56] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_g[55] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_g[54] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_g[53] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_g[52] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_g[51] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_g[50] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_g[49] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_g[48] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_g[47] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_g[46] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_g[45] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_g[44] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_g[43] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_g[42] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_g[41] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_g[40] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[61]=i_g[60] | i_p[60]&i_g[59] | i_p[60]&i_p[59]&i_g[58] | i_p[60]&i_p[59]&i_p[58]&i_g[57] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_g[56] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_g[55] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_g[54] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_g[53] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_g[52] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_g[51] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_g[50] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_g[49] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_g[48] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_g[47] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_g[46] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_g[45] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_g[44] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_g[43] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_g[42] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_g[41] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_g[40] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[62]=i_g[61] | i_p[61]&i_g[60] | i_p[61]&i_p[60]&i_g[59] | i_p[61]&i_p[60]&i_p[59]&i_g[58] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_g[57] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_g[56] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_g[55] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_g[54] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_g[53] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_g[52] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_g[51] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_g[50] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_g[49] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_g[48] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_g[47] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_g[46] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_g[45] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_g[44] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_g[43] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_g[42] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_g[41] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_g[40] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[63]=i_g[62] | i_p[62]&i_g[61] | i_p[62]&i_p[61]&i_g[60] | i_p[62]&i_p[61]&i_p[60]&i_g[59] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_g[58] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_g[57] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_g[56] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_g[55] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_g[54] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_g[53] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_g[52] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_g[51] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_g[50] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_g[49] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_g[48] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_g[47] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_g[46] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_g[45] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_g[44] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_g[43] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_g[42] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_g[41] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_g[40] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[64]=i_g[63] | i_p[63]&i_g[62] | i_p[63]&i_p[62]&i_g[61] | i_p[63]&i_p[62]&i_p[61]&i_g[60] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_g[59] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_g[58] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_g[57] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_g[56] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_g[55] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_g[54] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_g[53] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_g[52] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_g[51] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_g[50] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_g[49] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_g[48] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_g[47] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_g[46] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_g[45] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_g[44] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_g[43] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_g[42] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_g[41] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_g[40] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;

/*
wire c0_63=i_g[62] | i_p[62]&i_g[61] | i_p[62]&i_p[61]&i_g[60] | i_p[62]&i_p[61]&i_p[60]&i_g[59] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_g[58] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_g[57] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_g[56] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_g[55] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_g[54] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_g[53] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_g[52] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_g[51] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_g[50] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_g[49] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_g[48] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_g[47] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_g[46] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_g[45] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_g[44] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_g[43] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_g[42] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_g[41] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_g[40] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23]; 
wire c1_63=i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[63]=c0_63 | c1_63; // sublime 超过极限宽度了，字体都变灰色了。因此将信号分成两部分书写

wire c0_64=i_g[63] | i_p[63]&i_g[62] | i_p[63]&i_p[62]&i_g[61] | i_p[63]&i_p[62]&i_p[61]&i_g[60] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_g[59] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_g[58] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_g[57] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_g[56] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_g[55] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_g[54] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_g[53] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_g[52] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_g[51] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_g[50] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_g[49] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_g[48] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_g[47] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_g[46] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_g[45] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_g[44] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_g[43] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_g[42] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_g[41] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_g[40] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23]; 
wire c1_64=i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_p[ 0]&i_c;
assign o_c[64]=c0_64 | c1_64;


wire gm0=i_g[63] | i_p[63]&i_g[62] | i_p[63]&i_p[62]&i_g[61] | i_p[63]&i_p[62]&i_p[61]&i_g[60] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_g[59] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_g[58] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_g[57] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_g[56] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_g[55] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_g[54] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_g[53] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_g[52] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_g[51] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_g[50] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_g[49] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_g[48] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_g[47] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_g[46] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_g[45] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_g[44] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_g[43] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_g[42] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_g[41] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_g[40] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23]; 
wire gm1=i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0];
assign o_gm=gm0 | gm1;
*/
assign o_gm=i_g[63] | i_p[63]&i_g[62] | i_p[63]&i_p[62]&i_g[61] | i_p[63]&i_p[62]&i_p[61]&i_g[60] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_g[59] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_g[58] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_g[57] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_g[56] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_g[55] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_g[54] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_g[53] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_g[52] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_g[51] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_g[50] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_g[49] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_g[48] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_g[47] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_g[46] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_g[45] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_g[44] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_g[43] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_g[42] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_g[41] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_g[40] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_g[39] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_g[38] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_g[37] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_g[36] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_g[35] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_g[34] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_g[33] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_g[32] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_g[31] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_g[30] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_g[29] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_g[28] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_g[27] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_g[26] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_g[25] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_g[24] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_g[23] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_g[22] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_g[21] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_g[20] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_g[19] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_g[18] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_g[17] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_g[16] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_g[15] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_g[14] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_g[13] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_g[12] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_g[11] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_g[10] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_g[ 9] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_g[ 8] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_g[ 7] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_g[ 6] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_g[ 5] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_g[ 4] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_g[ 3] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_g[ 2] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_g[ 1] | i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[ 9]&i_p[ 8]&i_p[ 7]&i_p[ 6]&i_p[ 5]&i_p[ 4]&i_p[ 3]&i_p[ 2]&i_p[ 1]&i_g[ 0];
assign o_pm=i_p[63]&i_p[62]&i_p[61]&i_p[60]&i_p[59]&i_p[58]&i_p[57]&i_p[56]&i_p[55]&i_p[54]&i_p[53]&i_p[52]&i_p[51]&i_p[50]&i_p[49]&i_p[48]&i_p[47]&i_p[46]&i_p[45]&i_p[44]&i_p[43]&i_p[42]&i_p[41]&i_p[40]&i_p[39]&i_p[38]&i_p[37]&i_p[36]&i_p[35]&i_p[34]&i_p[33]&i_p[32]&i_p[31]&i_p[30]&i_p[29]&i_p[28]&i_p[27]&i_p[26]&i_p[25]&i_p[24]&i_p[23]&i_p[22]&i_p[21]&i_p[20]&i_p[19]&i_p[18]&i_p[17]&i_p[16]&i_p[15]&i_p[14]&i_p[13]&i_p[12]&i_p[11]&i_p[10]&i_p[9]&i_p[8]&i_p[7]&i_p[6]&i_p[5]&i_p[4]&i_p[3]&i_p[2]&i_p[1]&i_p[0];// propagater of MSB
endmodule
